// NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE
// This is an automatically generated file by stavros on Τετ 02 Μαρ 2022 07:35:18 μμ EET
//
// cmd:    swerv -snapshot=swerv-app -unset=assert_on -set=reset_vec=0x80000000 -set=fpga_optimize=1 
//

`include "common_defines.vh"
`undef ASSERT_ON
`undef TEC_RV_ICG
`define TEC_RV_ICG CKLNQD12BWP35P140
`define PHYSICAL 1
